`timescale 1ps/1ps
module testbench();
    reg clk;
    reg n_rst;
    reg [7:0] data;
    reg valid;

    wire [3:0] dtype;
    wire [4:0] op;
    wire [15:0] src1;
    wire [15:0] src2;
    wire done;

    decorder dut_decorder (
        .clk(clk),
        .n_rst(n_rst),
        .data(data),
        .valid(valid),
        .dtype(dtype),
        .op(op),
        .src1(src1),
        .src2(src2),
        .done(done)
    );

    always #5 clk = ~clk;
    initial begin
        clk = 1'b0;
        n_rst = 1'b0;
        #7 n_rst = 1'b1;
    end

    initial begin
        data = 8'h00;
        valid = 1'b0;
        #22;
        data = 8'h48;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//real start
        data = 8'h49;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//space
        data = 8'h20;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//type
        data = 8'h53;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//data1_space
        data = 8'h20;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//d1_1
        data = 8'h31;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//d1_7
        data = 8'h37;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//d1_4
        data = 8'h34;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//d1_9
        data = 8'h39;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//op sub
        data = 8'h2d;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//data_2 want 1248 d2_1
        data = 8'h31;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//d2_2
        data = 8'h32;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//d2_4
        data = 8'h34;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//d2_8
        data = 8'h38;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//equal state
        data = 8'h2b;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #40;
//equal = 3d
        data = 8'h3d;
        #10;
        valid = 1'b1;
        #10;
        valid = 1'b0;
        #100;

        $stop;
    end

endmodule