`timescale 1ps/1ps
module testbench();
    reg [31:0] A;
    reg [31:0] B;
    reg c_in;
    wire [31:0] sum;
    wire c_out;


    initial begin



        $stop
    end


endmodule